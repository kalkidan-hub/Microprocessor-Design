module fsm(clk,reset,x,y);
    input clk,reset,x;
    output y;
    
endmodule